// test bech for sin module
`timescale 1ns/1ns

module sinTB ();
  reg clk = 0;
  reg rst = 0;
  reg start = 0;
  reg [15:0] xBus;
  wire done;
  wire [17:0] rBus;

  sinTop sin(clk, rst, start, xBus, rBus, done);

  // generating clock behaviour
  always #5 clk <= ~clk;
  initial begin
    // Dump waveform data to a file.
    $dumpfile("sin_sim.vcd");
    $dumpvars(0, sinTB);

    // x = 0 rad => sin(x) = 0.0 rad
    #5;
    rst = 1;

    #5;
    #5;
    rst = 0;
    xBus = 0;
    start = 1;

    #5;
    #5;
    start = 0;

    #300;

    // x = 0.125 rad => sin(x) = 0.12467 rad
    #5;
    rst = 1;

    #5;
    #5;
    rst = 0;
    xBus = 16'h2000; // 0.125
    start = 1;

    #5;
    #5;
    start = 0;

    #300;

    // x = 0.25 rad => sin(x) = 0.24740 rad
    #5;
    rst = 1;

    #5;
    #5;
    rst = 0;
    xBus = 16'h4000; // 0.25
    start = 1;

    #5;
    #5;
    start = 0;

    #300;
    // x = 0.5 rad => sin(x) = 0.479425 rad
    #5;
    rst = 1;

    #5;
    #5;
    rst = 0;
    xBus = 16'h8000; // 0.5
    start = 1;

    #5;
    #5;
    start = 0;

    #300;
    // x = 1 rad => sin(x) = 0.84147 rad
    #5;
    rst = 1;

    #5;
    #5;
    rst = 0;
    xBus = 16'hFFFF; // 1 
    start = 1;

    #5;
    #5;
    start = 0;

    #300;

    // x = 1.5 rad => sin(1.5) ≈ 0.99749
    #5; rst = 1;
    #5; #5; rst = 0; xBus = 16'h18000; start = 1;
    #5; #5; start = 0;
    #300;

    // x = 2 rad => sin(2) ≈ 0.90929
    #5; rst = 1;
    #5; #5; rst = 0; xBus = 16'h20000; start = 1;
    #5; #5; start = 0;
    #300;

    // x = 2.5 rad => sin(2.5) ≈ 0.59847
    #5; rst = 1;
    #5; #5; rst = 0; xBus = 16'h28000; start = 1;
    #5; #5; start = 0;
    #300;

    // x = 3 rad => sin(3) ≈ 0.14112
    #5; rst = 1;
    #5; #5; rst = 0; xBus = 16'h30000; start = 1;
    #5; #5; start = 0;
    #300;

    // x = 3.5 rad => sin(3.5) ≈ -0.35078
    #5; rst = 1;
    #5; #5; rst = 0; xBus = 16'h38000; start = 1;
    #5; #5; start = 0;
    #300;

    $finish; 
  end

endmodule
